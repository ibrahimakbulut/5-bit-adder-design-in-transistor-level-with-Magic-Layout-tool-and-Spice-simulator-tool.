* SPICE3 file created from adder.ext - technology: scmos

.option scale=0.12u

M1000 xor2_0/nand2_1/a bin vdd xor2_0/nand2_0/w_n15_7# pmos w=18 l=2
+  ad=108 pd=48 as=2340 ps=1196
M1001 vdd bin xor2_0/nand2_1/a xor2_0/nand2_0/w_n15_7# pmos w=18 l=2
+  ad=0 pd=0 as=0 ps=0
M1002 xor2_0/nand2_0/a_n2_n7# bin gnd gnd nmos w=8 l=2
+  ad=32 pd=24 as=520 ps=338
M1003 xor2_0/nand2_1/a bin xor2_0/nand2_0/a_n2_n7# gnd nmos w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1004 xor2_0/nand2_4/a xor2_0/nand2_1/a vdd xor2_0/nand2_1/w_n15_7# pmos w=18 l=2
+  ad=108 pd=48 as=0 ps=0
M1005 vdd ain xor2_0/nand2_4/a xor2_0/nand2_1/w_n15_7# pmos w=18 l=2
+  ad=0 pd=0 as=0 ps=0
M1006 xor2_0/nand2_1/a_n2_n7# xor2_0/nand2_1/a gnd gnd nmos w=8 l=2
+  ad=32 pd=24 as=0 ps=0
M1007 xor2_0/nand2_4/a ain xor2_0/nand2_1/a_n2_n7# gnd nmos w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1008 xor2_0/nand2_3/a ain vdd xor2_0/nand2_2/w_n15_7# pmos w=18 l=2
+  ad=108 pd=48 as=0 ps=0
M1009 vdd ain xor2_0/nand2_3/a xor2_0/nand2_2/w_n15_7# pmos w=18 l=2
+  ad=0 pd=0 as=0 ps=0
M1010 xor2_0/nand2_2/a_n2_n7# ain gnd gnd nmos w=8 l=2
+  ad=32 pd=24 as=0 ps=0
M1011 xor2_0/nand2_3/a ain xor2_0/nand2_2/a_n2_n7# gnd nmos w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1012 xor2_0/nand2_4/b xor2_0/nand2_3/a vdd xor2_0/nand2_3/w_n15_7# pmos w=18 l=2
+  ad=108 pd=48 as=0 ps=0
M1013 vdd bin xor2_0/nand2_4/b xor2_0/nand2_3/w_n15_7# pmos w=18 l=2
+  ad=0 pd=0 as=0 ps=0
M1014 xor2_0/nand2_3/a_n2_n7# xor2_0/nand2_3/a gnd gnd nmos w=8 l=2
+  ad=32 pd=24 as=0 ps=0
M1015 xor2_0/nand2_4/b bin xor2_0/nand2_3/a_n2_n7# gnd nmos w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1016 nand2_0/a xor2_0/nand2_4/a vdd xor2_0/nand2_4/w_n15_7# pmos w=18 l=2
+  ad=108 pd=48 as=0 ps=0
M1017 vdd xor2_0/nand2_4/b nand2_0/a xor2_0/nand2_4/w_n15_7# pmos w=18 l=2
+  ad=0 pd=0 as=0 ps=0
M1018 xor2_0/nand2_4/a_n2_n7# xor2_0/nand2_4/a gnd gnd nmos w=8 l=2
+  ad=32 pd=24 as=0 ps=0
M1019 nand2_0/a xor2_0/nand2_4/b xor2_0/nand2_4/a_n2_n7# gnd nmos w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1020 xor2_1/nand2_1/a nand2_0/a vdd xor2_1/nand2_0/w_n15_7# pmos w=18 l=2
+  ad=108 pd=48 as=0 ps=0
M1021 vdd nand2_0/a xor2_1/nand2_1/a xor2_1/nand2_0/w_n15_7# pmos w=18 l=2
+  ad=0 pd=0 as=0 ps=0
M1022 xor2_1/nand2_0/a_n2_n7# nand2_0/a gnd gnd nmos w=8 l=2
+  ad=32 pd=24 as=0 ps=0
M1023 xor2_1/nand2_1/a nand2_0/a xor2_1/nand2_0/a_n2_n7# gnd nmos w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1024 xor2_1/nand2_4/a xor2_1/nand2_1/a vdd xor2_1/nand2_1/w_n15_7# pmos w=18 l=2
+  ad=108 pd=48 as=0 ps=0
M1025 vdd cin xor2_1/nand2_4/a xor2_1/nand2_1/w_n15_7# pmos w=18 l=2
+  ad=0 pd=0 as=0 ps=0
M1026 xor2_1/nand2_1/a_n2_n7# xor2_1/nand2_1/a gnd gnd nmos w=8 l=2
+  ad=32 pd=24 as=0 ps=0
M1027 xor2_1/nand2_4/a cin xor2_1/nand2_1/a_n2_n7# gnd nmos w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1028 xor2_1/nand2_3/a cin vdd xor2_1/nand2_2/w_n15_7# pmos w=18 l=2
+  ad=108 pd=48 as=0 ps=0
M1029 vdd cin xor2_1/nand2_3/a xor2_1/nand2_2/w_n15_7# pmos w=18 l=2
+  ad=0 pd=0 as=0 ps=0
M1030 xor2_1/nand2_2/a_n2_n7# cin gnd gnd nmos w=8 l=2
+  ad=32 pd=24 as=0 ps=0
M1031 xor2_1/nand2_3/a cin xor2_1/nand2_2/a_n2_n7# gnd nmos w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1032 xor2_1/nand2_4/b xor2_1/nand2_3/a vdd xor2_1/nand2_3/w_n15_7# pmos w=18 l=2
+  ad=108 pd=48 as=0 ps=0
M1033 vdd nand2_0/a xor2_1/nand2_4/b xor2_1/nand2_3/w_n15_7# pmos w=18 l=2
+  ad=0 pd=0 as=0 ps=0
M1034 xor2_1/nand2_3/a_n2_n7# xor2_1/nand2_3/a gnd gnd nmos w=8 l=2
+  ad=32 pd=24 as=0 ps=0
M1035 xor2_1/nand2_4/b nand2_0/a xor2_1/nand2_3/a_n2_n7# gnd nmos w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1036 sum xor2_1/nand2_4/a vdd xor2_1/nand2_4/w_n15_7# pmos w=18 l=2
+  ad=108 pd=48 as=0 ps=0
M1037 vdd xor2_1/nand2_4/b sum xor2_1/nand2_4/w_n15_7# pmos w=18 l=2
+  ad=0 pd=0 as=0 ps=0
M1038 xor2_1/nand2_4/a_n2_n7# xor2_1/nand2_4/a gnd gnd nmos w=8 l=2
+  ad=32 pd=24 as=0 ps=0
M1039 sum xor2_1/nand2_4/b xor2_1/nand2_4/a_n2_n7# gnd nmos w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1040 nand2_2/b nand2_0/a vdd nand2_0/w_n15_7# pmos w=18 l=2
+  ad=108 pd=48 as=0 ps=0
M1041 vdd cin nand2_2/b nand2_0/w_n15_7# pmos w=18 l=2
+  ad=0 pd=0 as=0 ps=0
M1042 nand2_0/a_n2_n7# nand2_0/a gnd gnd nmos w=8 l=2
+  ad=32 pd=24 as=0 ps=0
M1043 nand2_2/b cin nand2_0/a_n2_n7# gnd nmos w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1044 nand2_2/a bin vdd nand2_1/w_n15_7# pmos w=18 l=2
+  ad=108 pd=48 as=0 ps=0
M1045 vdd ain nand2_2/a nand2_1/w_n15_7# pmos w=18 l=2
+  ad=0 pd=0 as=0 ps=0
M1046 nand2_1/a_n2_n7# bin gnd gnd nmos w=8 l=2
+  ad=32 pd=24 as=0 ps=0
M1047 nand2_2/a ain nand2_1/a_n2_n7# gnd nmos w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1048 cout nand2_2/a vdd nand2_2/w_n15_7# pmos w=18 l=2
+  ad=108 pd=48 as=0 ps=0
M1049 vdd nand2_2/b cout nand2_2/w_n15_7# pmos w=18 l=2
+  ad=0 pd=0 as=0 ps=0
M1050 nand2_2/a_n2_n7# nand2_2/a gnd gnd nmos w=8 l=2
+  ad=32 pd=24 as=0 ps=0
M1051 cout nand2_2/b nand2_2/a_n2_n7# gnd nmos w=8 l=2
+  ad=40 pd=26 as=0 ps=0
C0 xor2_1/nand2_4/w_n15_7# xor2_1/nand2_4/a 0.11fF
C1 cout cin 0.01fF
C2 nand2_2/a nand2_2/w_n15_7# 0.14fF
C3 nand2_0/w_n15_7# cout 0.03fF
C4 xor2_1/nand2_3/w_n15_7# xor2_1/nand2_3/a 0.14fF
C5 xor2_1/nand2_2/w_n15_7# xor2_1/nand2_3/a 0.06fF
C6 xor2_0/nand2_1/a_n2_n7# vdd 0.01fF
C7 vdd nand2_2/b 0.45fF
C8 bin xor2_0/nand2_3/a 0.09fF
C9 xor2_1/nand2_1/w_n15_7# xor2_1/nand2_4/a 0.06fF
C10 cout vdd 0.58fF
C11 xor2_0/nand2_4/w_n15_7# xor2_0/nand2_4/a 0.11fF
C12 xor2_0/nand2_0/w_n15_7# bin 0.24fF
C13 xor2_1/nand2_1/w_n15_7# xor2_1/nand2_1/a 0.14fF
C14 xor2_0/nand2_3/a gnd 0.08fF
C15 xor2_0/nand2_1/a xor2_0/nand2_0/w_n15_7# 0.06fF
C16 gnd nand2_2/a 0.08fF
C17 xor2_1/nand2_1/a xor2_1/nand2_4/a 0.05fF
C18 xor2_0/nand2_3/w_n15_7# xor2_0/nand2_3/a 0.14fF
C19 gnd xor2_1/nand2_4/w_n15_7# 0.01fF
C20 vdd xor2_1/nand2_1/a_n2_n7# 0.01fF
C21 ain xor2_0/nand2_3/a 0.03fF
C22 ain nand2_2/a 0.03fF
C23 xor2_1/nand2_4/w_n15_7# xor2_1/nand2_4/b 0.11fF
C24 xor2_0/nand2_4/b xor2_0/nand2_3/a 0.05fF
C25 nand2_0/a xor2_1/nand2_3/w_n15_7# 0.11fF
C26 xor2_1/nand2_3/w_n15_7# xor2_1/nand2_4/b 0.06fF
C27 sum gnd 0.04fF
C28 xor2_0/nand2_1/w_n15_7# xor2_0/nand2_1/a 0.14fF
C29 sum xor2_1/nand2_4/b 0.03fF
C30 gnd xor2_1/nand2_4/a 0.04fF
C31 cin xor2_1/nand2_2/w_n15_7# 0.24fF
C32 gnd xor2_1/nand2_3/a 0.08fF
C33 xor2_1/nand2_4/a xor2_1/nand2_4/b 0.09fF
C34 nand2_0/a xor2_1/nand2_3/a 0.09fF
C35 gnd xor2_1/nand2_1/a 0.08fF
C36 xor2_0/nand2_3/a vdd 0.49fF
C37 xor2_1/nand2_3/a xor2_1/nand2_4/b 0.05fF
C38 nand2_2/a vdd 0.49fF
C39 xor2_1/nand2_1/w_n15_7# cin 0.13fF
C40 xor2_0/nand2_1/a bin 0.03fF
C41 nand2_0/a xor2_1/nand2_1/a 0.03fF
C42 vdd xor2_1/nand2_4/w_n15_7# 0.18fF
C43 cin xor2_1/nand2_4/a 0.03fF
C44 xor2_0/nand2_1/w_n15_7# ain 0.13fF
C45 xor2_0/nand2_0/w_n15_7# vdd 0.17fF
C46 vdd xor2_1/nand2_3/w_n15_7# 0.18fF
C47 cin xor2_1/nand2_3/a 0.03fF
C48 bin gnd 0.94fF
C49 vdd xor2_1/nand2_2/w_n15_7# 0.17fF
C50 xor2_0/nand2_1/a gnd 0.08fF
C51 cout nand2_2/b 0.13fF
C52 xor2_1/nand2_1/a cin 0.09fF
C53 bin xor2_0/nand2_3/w_n15_7# 0.11fF
C54 sum vdd 0.45fF
C55 xor2_1/nand2_1/w_n15_7# vdd 0.17fF
C56 ain bin 1.17fF
C57 vdd xor2_1/nand2_4/a 0.72fF
C58 bin xor2_0/nand2_4/b 0.03fF
C59 xor2_0/nand2_1/a ain 0.09fF
C60 gnd nand2_0/a 1.04fF
C61 vdd xor2_1/nand2_3/a 0.49fF
C62 gnd xor2_1/nand2_4/b 0.36fF
C63 xor2_0/nand2_1/w_n15_7# vdd 0.17fF
C64 xor2_0/nand2_2/w_n15_7# xor2_0/nand2_3/a 0.06fF
C65 vdd nand2_2/w_n15_7# 0.17fF
C66 xor2_1/nand2_0/w_n15_7# xor2_1/nand2_1/a 0.06fF
C67 ain gnd 0.10fF
C68 nand2_0/a xor2_1/nand2_4/b 0.03fF
C69 xor2_1/nand2_1/a vdd 0.54fF
C70 nand2_1/w_n15_7# nand2_2/a 0.06fF
C71 xor2_0/nand2_4/b gnd 0.36fF
C72 gnd cin 0.10fF
C73 xor2_0/nand2_4/b nand2_0/a 0.03fF
C74 xor2_0/nand2_3/w_n15_7# xor2_0/nand2_4/b 0.06fF
C75 nand2_0/a cin 1.09fF
C76 bin vdd 0.72fF
C77 nand2_0/w_n15_7# nand2_0/a 0.11fF
C78 xor2_0/nand2_1/a vdd 0.54fF
C79 nand2_2/a nand2_2/b 0.09fF
C80 nand2_0/w_n15_7# cin 0.13fF
C81 gnd vdd 0.31fF
C82 xor2_1/nand2_0/w_n15_7# nand2_0/a 0.24fF
C83 nand2_0/a vdd 1.01fF
C84 xor2_0/nand2_3/w_n15_7# vdd 0.18fF
C85 vdd xor2_1/nand2_4/b 0.45fF
C86 nand2_2/a cout 0.07fF
C87 ain vdd 0.43fF
C88 xor2_0/nand2_4/b vdd 0.45fF
C89 xor2_0/nand2_1/w_n15_7# xor2_0/nand2_4/a 0.06fF
C90 cin vdd 0.55fF
C91 nand2_0/w_n15_7# vdd 0.16fF
C92 gnd xor2_0/nand2_4/w_n15_7# 0.01fF
C93 nand2_1/w_n15_7# bin 0.11fF
C94 xor2_0/nand2_4/w_n15_7# nand2_0/a 0.06fF
C95 nand2_2/w_n15_7# nand2_2/b 0.11fF
C96 xor2_1/nand2_0/w_n15_7# vdd 0.17fF
C97 xor2_0/nand2_1/a xor2_0/nand2_4/a 0.05fF
C98 xor2_0/nand2_4/b xor2_0/nand2_4/w_n15_7# 0.11fF
C99 cout nand2_2/w_n15_7# 0.06fF
C100 gnd xor2_0/nand2_4/a 0.04fF
C101 ain xor2_0/nand2_2/w_n15_7# 0.24fF
C102 ain nand2_1/w_n15_7# 0.13fF
C103 ain xor2_0/nand2_4/a 0.03fF
C104 gnd nand2_2/b 0.37fF
C105 xor2_0/nand2_4/b xor2_0/nand2_4/a 0.09fF
C106 xor2_0/nand2_4/w_n15_7# vdd 0.18fF
C107 gnd cout 0.30fF
C108 xor2_0/nand2_2/w_n15_7# vdd 0.17fF
C109 nand2_0/a cout 0.01fF
C110 nand2_1/w_n15_7# vdd 0.17fF
C111 cin nand2_2/b 0.03fF
C112 sum xor2_1/nand2_4/w_n15_7# 0.06fF
C113 nand2_0/w_n15_7# nand2_2/b 0.06fF
C114 xor2_0/nand2_4/a vdd 0.72fF
C115 cout gnd 0.56fF
C116 nand2_2/a gnd 0.40fF
C117 nand2_2/w_n15_7# gnd 0.87fF
C118 nand2_1/w_n15_7# gnd 0.87fF
C119 nand2_2/b gnd 0.29fF
C120 nand2_0/w_n15_7# gnd 0.87fF
C121 gnd gnd 5.00fF
C122 sum gnd 0.12fF
C123 xor2_1/nand2_4/b gnd 0.45fF
C124 xor2_1/nand2_4/w_n15_7# gnd 0.87fF
C125 xor2_1/nand2_3/a gnd 0.34fF
C126 xor2_1/nand2_3/w_n15_7# gnd 0.87fF
C127 xor2_1/nand2_2/w_n15_7# gnd 0.87fF
C128 vdd gnd 3.02fF
C129 cin gnd 1.65fF
C130 xor2_1/nand2_1/a gnd 0.06fF
C131 xor2_1/nand2_1/w_n15_7# gnd 0.87fF
C132 nand2_0/a gnd 1.38fF
C133 xor2_1/nand2_0/w_n15_7# gnd 0.87fF
C134 xor2_0/nand2_4/b gnd 0.45fF
C135 xor2_0/nand2_4/w_n15_7# gnd 0.87fF
C136 xor2_0/nand2_3/a gnd 0.34fF
C137 xor2_0/nand2_3/w_n15_7# gnd 0.87fF
C138 xor2_0/nand2_2/w_n15_7# gnd 0.87fF
C139 ain gnd 1.73fF
C140 xor2_0/nand2_1/a gnd 0.06fF
C141 xor2_0/nand2_1/w_n15_7# gnd 0.87fF
C142 bin gnd 1.36fF
C143 xor2_0/nand2_0/w_n15_7# gnd 0.87fF


* INDEPENDANT VOLTAGE SOURCE
*
*Vname +NODE -NODE VALUE
*----- ----- ----- -----
VCC    vdd     gnd     DC=2.5
Vcin0  cin     gnd     DC=0

* The following two lines are for TRANSIENT analysis
*
*Vname +Node -Node Option T1  V1   T2  V2   T3   V3    T4  V4  T5   V5 
*----- ----- ----- ------ --  --   --  --   ---- --    --  --  ---- -- 
*V1     cin     gnd    PWL(   0N   0  0.1N  0  16N  0    16.1N 2.5   32N  2.5 32.1N 0) 
V2     ain     gnd    PWL(   0N   0  0.1N  0  8N  0    8.1N 2.5   16N  2.5 16.1N 0      24N  0    24.1N 2.5   32N  2.5 32.1N 0) 
V3     bin     gnd    PWL(   0N   0  0.1N  0  4N  0    4.1N 2.5   8N  2.5 8.1N 0      12N  0    12.1N 2.5   16N  2.5 16.1N 0    20N   0    20.1N  2.5    24N 2.5   24.1N  0 28N 0      28.1N  2.5    32N  2.5 32.1N 0) 


*     TSTEP TSTOP
*     ----- -----
.TRAN 0.1N  35N

* TEMPERATURE and OPTIONS SETTING

.OPTIONS TEMP=25 reltol = 1e-6

*MODELS

.include tsmc_cmos025

.END